version https://git-lfs.github.com/spec/v1
oid sha256:25f901f7169ad06685698d21ddefd322a5134c272edebbd39a4f894ec97e8658
size 1120
